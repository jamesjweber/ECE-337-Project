module tb_AES_block();

endmodule

module slave_read (

);

endmodule // slave_read

module()


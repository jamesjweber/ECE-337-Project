// 337 TA Provided Lab 2 Testbench
// This code serves as a starer test bench for the synchronizer design
// STUDENT: Replace this message and the above header section with an
// appropriate header based on your other code files

// 0.5um D-FlipFlop Timing Data Estimates:
// Data Propagation delay (clk->Q): 670ps
// Setup time for data relative to clock: 190ps
// Hold time for data relative to clock: 10ps

`timescale 1ns / 10ps

module tb_encryption_block();

	// Define local parameters used by the test bench
	localparam	CLK_PERIOD		= 5;
	//localparam	FF_SETUP_TIME	= 0.190;
	//localparam	FF_HOLD_TIME	= 0.100;
	//localparam	CHECK_DELAY 	= (CLK_PERIOD - FF_SETUP_TIME); // Check right before the setup time starts
	
	//localparam	RESET_OUTPUT_VALUE	= 1'b1;
	
	// Declare DUT portmap signals
	reg tb_clk;
	reg tb_rst;
	reg tb_keyLock;
	reg tb_go;
	reg tb_done;
	reg [2:0] tb_keySelect;
	reg [2:0] tb_encSelect;
	reg [4:0] tb_count;
	reg [127:0] tb_keyIn;
	reg [127:0] tb_nonceIn;
	reg [127:0] tb_pText;
	reg [127:0] tb_encText;
	
	// Declare test bench signals
	//integer tb_test_num;
	//string tb_test_case;
	//integer tb_stream_test_num;
	
	// Clock generation block
	always
	begin
		tb_clk = 1'b0;
		#(CLK_PERIOD/3.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD/3.0);
	end
	
	// DUT Port map
	encryption_block DUT(.clk(tb_clk), .rst(tb_rst), .keyLock(tb_keyLock), .fsmGo(tb_go), .done(tb_done), .count(tb_count), .keySelect(tb_keySelect), .encSelect(tb_encSelect), .keyIn(tb_keyIn), .nonceIn(tb_nonceIn), .pText(tb_pText), .encText(tb_encText));
	// Test bench main process
	initial
	begin
		tb_count = 0;
		tb_rst = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyIn = 127'b0;
		tb_nonceIn = 127'b0;
		tb_keySelect = 3'b011;
		tb_encSelect = 3'b000;
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_rst = 1'b0;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_go = 1;
		tb_keySelect = tb_keySelect - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_keySelect = tb_keySelect - 1;
		tb_encSelect = tb_encSelect + 1;
		tb_count = tb_count + 1;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_go = 0;
		tb_pText = 128'hFFFF;
		@(posedge tb_clk);	
		tb_pText = 128'hF00F;	
		@(posedge tb_clk);
		tb_pText = 128'h0FF0;
		@(posedge tb_clk);
		tb_pText = 128'h0FF0;
		@(posedge tb_clk);

	end
endmodule
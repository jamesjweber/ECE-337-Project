module tb_ahb_lite_slave_interface();

endmodule

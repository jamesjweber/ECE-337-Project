`timescale 1ns / 10ps

module tb_key_block();

	localparam CLK_PERIOD = 5;

	// Declare DUT portmap signals
	reg tb_clk;
	reg tb_rst;
	reg tb_keyLock;
	reg [2:0] tb_select;
	reg [127:0] tb_in;
	reg [127:0] tb_roundKey;
	reg [127:0] tb_froundKey;
	
	// Clock generation block
	always
	begin
		tb_clk = 1'b0;
		#(CLK_PERIOD/3.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD/3.0);
	end
	
	// DUT Port map
	key_block DUT(.clk(tb_clk), .rst(tb_rst), .keyLock(tb_keyLock), .select(tb_select), .in(tb_in), .roundKey(tb_roundKey), .froundKey(tb_froundKey));

	// Test bench main process
	initial
	begin
		tb_rst = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_in = 128'h0123456789ABCDEF0123456789ABCDEF;
		tb_select = 6'b011;
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_rst = 1'b0;
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
		tb_select = tb_select - 1; 	
		@(posedge tb_clk);		
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_keyLock = 1;
		@(posedge tb_clk);
		tb_keyLock = 0;
	end
endmodule

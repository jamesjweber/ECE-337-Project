module s_box
(
	input wire [2:0] sel,
	input wire [127:0] inData,
	output reg [127:0] outData
);

	reg [0:15] S0 = {4'd3, 4'd8, 4'd15, 4'd1, 4'd10, 4'd6, 4'd5, 4'd11, 4'd14, 4'd13, 4'd4, 4'd2, 4'd7, 4'd0, 4'd9, 4'd12};
	reg [0:15] S1 = {4'd15, 4'd12, 4'd2, 4'd7, 4'd9, 4'd0, 4'd5, 4'd10, 4'd1, 4'd11, 4'd14, 4'd8, 4'd6, 4'd13, 4'd3, 4'd4};
	reg [0:15] S2 = {4'd8, 4'd6, 4'd7, 4'd9, 4'd3, 4'd12, 4'd10, 4'd15, 4'd13, 4'd1, 4'd14, 4'd4, 4'd0, 4'd11, 4'd5, 4'd2};
	reg [0:15] S3 = {4'd0, 4'd15, 4'd11, 4'd8, 4'd12, 4'd9, 4'd6, 4'd3, 4'd13, 4'd1, 4'd2, 4'd4, 4'd10, 4'd7, 4'd5, 4'd14};
	reg [0:15] S4 = {4'd1, 4'd15, 4'd8, 4'd3, 4'd12, 4'd0, 4'd11, 4'd6, 4'd2, 4'd5, 4'd4, 4'd10, 4'd9, 4'd14, 4'd7, 4'd13};
	reg [0:15] S5 = {4'd15, 4'd5, 4'd2, 4'd11, 4'd4, 4'd10, 4'd9, 4'd12, 4'd0, 4'd3, 4'd14, 4'd8, 4'd13, 4'd6, 4'd7, 4'd1};
	reg [0:15] S6 = {4'd7, 4'd2, 4'd12, 4'd5, 4'd8, 4'd4, 4'd6, 4'd11, 4'd14, 4'd9, 4'd1, 4'd15, 4'd13, 4'd3, 4'd10, 4'd0};
	reg [0:15] S7 = {4'd1, 4'd13, 4'd15, 4'd0, 4'd14, 4'd8, 4'd2, 4'd11, 4'd7, 4'd4, 4'd12, 4'd10, 4'd9, 4'd3, 4'd5, 4'd6};

	reg [0:15] sBlocks [0:7] = {S0, S1, S2, S3, S4, S5, S6, S7};

	integer i;
	always_comb
	begin
		for(i = 3; i < 128; i += 4)
			outData[i-:3] = sBlocks[sel][inData[i-:3]];
	end

endmodule